// nios_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clk_clk,                //             clk.clk
		output wire [9:0]  doodle_x_export,        //        doodle_x.export
		output wire [9:0]  doodle_y_export,        //        doodle_y.export
		output wire [9:0]  floor1_x_export,        //        floor1_x.export
		output wire [9:0]  floor1_y_export,        //        floor1_y.export
		output wire [9:0]  floor2_x_export,        //        floor2_x.export
		output wire [9:0]  floor2_y_export,        //        floor2_y.export
		output wire [9:0]  floor3_x_export,        //        floor3_x.export
		output wire [9:0]  floor3_y_export,        //        floor3_y.export
		output wire [9:0]  floor4_x_export,        //        floor4_x.export
		output wire [9:0]  floor4_y_export,        //        floor4_y.export
		output wire [9:0]  floor5_x_export,        //        floor5_x.export
		output wire [9:0]  floor5_y_export,        //        floor5_y.export
		output wire [9:0]  floor6_x_export,        //        floor6_x.export
		output wire [9:0]  floor6_y_export,        //        floor6_y.export
		output wire [9:0]  floor7_x_export,        //        floor7_x.export
		output wire [9:0]  floor7_y_export,        //        floor7_y.export
		output wire [9:0]  floor8_x_export,        //        floor8_x.export
		output wire [9:0]  floor8_y_export,        //        floor8_y.export
		output wire [7:0]  keycode_export,         //         keycode.export
		output wire [1:0]  otg_hpi_address_export, // otg_hpi_address.export
		output wire        otg_hpi_cs_export,      //      otg_hpi_cs.export
		input  wire [15:0] otg_hpi_data_in_port,   //    otg_hpi_data.in_port
		output wire [15:0] otg_hpi_data_out_port,  //                .out_port
		output wire        otg_hpi_r_export,       //       otg_hpi_r.export
		output wire        otg_hpi_reset_export,   //   otg_hpi_reset.export
		output wire        otg_hpi_w_export,       //       otg_hpi_w.export
		input  wire        reset_reset_n,          //           reset.reset_n
		output wire [15:0] score_export,           //           score.export
		output wire        sdram_clk_clk,          //       sdram_clk.clk
		output wire [12:0] sdram_wire_addr,        //      sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,          //                .ba
		output wire        sdram_wire_cas_n,       //                .cas_n
		output wire        sdram_wire_cke,         //                .cke
		output wire        sdram_wire_cs_n,        //                .cs_n
		inout  wire [31:0] sdram_wire_dq,          //                .dq
		output wire [3:0]  sdram_wire_dqm,         //                .dqm
		output wire        sdram_wire_ras_n,       //                .ras_n
		output wire        sdram_wire_we_n         //                .we_n
	);

	wire         sdram_pll_c0_clk;                                             // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_002:clk, sdram:clk]
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [28:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [28:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;        // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;         // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;               // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;                // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                   // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                  // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;              // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                        // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                          // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                       // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                           // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                              // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                        // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                     // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                             // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                         // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire   [7:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [18:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire   [7:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_doodle_x_s1_chipselect;                     // mm_interconnect_0:doodle_x_s1_chipselect -> doodle_x:chipselect
	wire  [31:0] mm_interconnect_0_doodle_x_s1_readdata;                       // doodle_x:readdata -> mm_interconnect_0:doodle_x_s1_readdata
	wire   [1:0] mm_interconnect_0_doodle_x_s1_address;                        // mm_interconnect_0:doodle_x_s1_address -> doodle_x:address
	wire         mm_interconnect_0_doodle_x_s1_write;                          // mm_interconnect_0:doodle_x_s1_write -> doodle_x:write_n
	wire  [31:0] mm_interconnect_0_doodle_x_s1_writedata;                      // mm_interconnect_0:doodle_x_s1_writedata -> doodle_x:writedata
	wire         mm_interconnect_0_doodle_y_s1_chipselect;                     // mm_interconnect_0:doodle_y_s1_chipselect -> doodle_y:chipselect
	wire  [31:0] mm_interconnect_0_doodle_y_s1_readdata;                       // doodle_y:readdata -> mm_interconnect_0:doodle_y_s1_readdata
	wire   [1:0] mm_interconnect_0_doodle_y_s1_address;                        // mm_interconnect_0:doodle_y_s1_address -> doodle_y:address
	wire         mm_interconnect_0_doodle_y_s1_write;                          // mm_interconnect_0:doodle_y_s1_write -> doodle_y:write_n
	wire  [31:0] mm_interconnect_0_doodle_y_s1_writedata;                      // mm_interconnect_0:doodle_y_s1_writedata -> doodle_y:writedata
	wire         mm_interconnect_0_floor1_x_s1_chipselect;                     // mm_interconnect_0:floor1_x_s1_chipselect -> floor1_x:chipselect
	wire  [31:0] mm_interconnect_0_floor1_x_s1_readdata;                       // floor1_x:readdata -> mm_interconnect_0:floor1_x_s1_readdata
	wire   [1:0] mm_interconnect_0_floor1_x_s1_address;                        // mm_interconnect_0:floor1_x_s1_address -> floor1_x:address
	wire         mm_interconnect_0_floor1_x_s1_write;                          // mm_interconnect_0:floor1_x_s1_write -> floor1_x:write_n
	wire  [31:0] mm_interconnect_0_floor1_x_s1_writedata;                      // mm_interconnect_0:floor1_x_s1_writedata -> floor1_x:writedata
	wire         mm_interconnect_0_floor1_y_s1_chipselect;                     // mm_interconnect_0:floor1_y_s1_chipselect -> floor1_y:chipselect
	wire  [31:0] mm_interconnect_0_floor1_y_s1_readdata;                       // floor1_y:readdata -> mm_interconnect_0:floor1_y_s1_readdata
	wire   [1:0] mm_interconnect_0_floor1_y_s1_address;                        // mm_interconnect_0:floor1_y_s1_address -> floor1_y:address
	wire         mm_interconnect_0_floor1_y_s1_write;                          // mm_interconnect_0:floor1_y_s1_write -> floor1_y:write_n
	wire  [31:0] mm_interconnect_0_floor1_y_s1_writedata;                      // mm_interconnect_0:floor1_y_s1_writedata -> floor1_y:writedata
	wire         mm_interconnect_0_keycode_s1_chipselect;                      // mm_interconnect_0:keycode_s1_chipselect -> keycode:chipselect
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                        // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                         // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire         mm_interconnect_0_keycode_s1_write;                           // mm_interconnect_0:keycode_s1_write -> keycode:write_n
	wire  [31:0] mm_interconnect_0_keycode_s1_writedata;                       // mm_interconnect_0:keycode_s1_writedata -> keycode:writedata
	wire         mm_interconnect_0_otg_hpi_address_s1_chipselect;              // mm_interconnect_0:otg_hpi_address_s1_chipselect -> otg_hpi_address:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_readdata;                // otg_hpi_address:readdata -> mm_interconnect_0:otg_hpi_address_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_address_s1_address;                 // mm_interconnect_0:otg_hpi_address_s1_address -> otg_hpi_address:address
	wire         mm_interconnect_0_otg_hpi_address_s1_write;                   // mm_interconnect_0:otg_hpi_address_s1_write -> otg_hpi_address:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_writedata;               // mm_interconnect_0:otg_hpi_address_s1_writedata -> otg_hpi_address:writedata
	wire         mm_interconnect_0_otg_hpi_data_s1_chipselect;                 // mm_interconnect_0:otg_hpi_data_s1_chipselect -> otg_hpi_data:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_readdata;                   // otg_hpi_data:readdata -> mm_interconnect_0:otg_hpi_data_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_data_s1_address;                    // mm_interconnect_0:otg_hpi_data_s1_address -> otg_hpi_data:address
	wire         mm_interconnect_0_otg_hpi_data_s1_write;                      // mm_interconnect_0:otg_hpi_data_s1_write -> otg_hpi_data:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_writedata;                  // mm_interconnect_0:otg_hpi_data_s1_writedata -> otg_hpi_data:writedata
	wire         mm_interconnect_0_otg_hpi_r_s1_chipselect;                    // mm_interconnect_0:otg_hpi_r_s1_chipselect -> otg_hpi_r:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_readdata;                      // otg_hpi_r:readdata -> mm_interconnect_0:otg_hpi_r_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_r_s1_address;                       // mm_interconnect_0:otg_hpi_r_s1_address -> otg_hpi_r:address
	wire         mm_interconnect_0_otg_hpi_r_s1_write;                         // mm_interconnect_0:otg_hpi_r_s1_write -> otg_hpi_r:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_writedata;                     // mm_interconnect_0:otg_hpi_r_s1_writedata -> otg_hpi_r:writedata
	wire         mm_interconnect_0_otg_hpi_cs_s1_chipselect;                   // mm_interconnect_0:otg_hpi_cs_s1_chipselect -> otg_hpi_cs:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_readdata;                     // otg_hpi_cs:readdata -> mm_interconnect_0:otg_hpi_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_cs_s1_address;                      // mm_interconnect_0:otg_hpi_cs_s1_address -> otg_hpi_cs:address
	wire         mm_interconnect_0_otg_hpi_cs_s1_write;                        // mm_interconnect_0:otg_hpi_cs_s1_write -> otg_hpi_cs:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_writedata;                    // mm_interconnect_0:otg_hpi_cs_s1_writedata -> otg_hpi_cs:writedata
	wire         mm_interconnect_0_otg_hpi_w_s1_chipselect;                    // mm_interconnect_0:otg_hpi_w_s1_chipselect -> otg_hpi_w:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_readdata;                      // otg_hpi_w:readdata -> mm_interconnect_0:otg_hpi_w_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_w_s1_address;                       // mm_interconnect_0:otg_hpi_w_s1_address -> otg_hpi_w:address
	wire         mm_interconnect_0_otg_hpi_w_s1_write;                         // mm_interconnect_0:otg_hpi_w_s1_write -> otg_hpi_w:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_writedata;                     // mm_interconnect_0:otg_hpi_w_s1_writedata -> otg_hpi_w:writedata
	wire         mm_interconnect_0_otg_hpi_reset_s1_chipselect;                // mm_interconnect_0:otg_hpi_reset_s1_chipselect -> otg_hpi_reset:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_readdata;                  // otg_hpi_reset:readdata -> mm_interconnect_0:otg_hpi_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_reset_s1_address;                   // mm_interconnect_0:otg_hpi_reset_s1_address -> otg_hpi_reset:address
	wire         mm_interconnect_0_otg_hpi_reset_s1_write;                     // mm_interconnect_0:otg_hpi_reset_s1_write -> otg_hpi_reset:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_writedata;                 // mm_interconnect_0:otg_hpi_reset_s1_writedata -> otg_hpi_reset:writedata
	wire         mm_interconnect_0_floor2_x_s1_chipselect;                     // mm_interconnect_0:floor2_x_s1_chipselect -> floor2_x:chipselect
	wire  [31:0] mm_interconnect_0_floor2_x_s1_readdata;                       // floor2_x:readdata -> mm_interconnect_0:floor2_x_s1_readdata
	wire   [1:0] mm_interconnect_0_floor2_x_s1_address;                        // mm_interconnect_0:floor2_x_s1_address -> floor2_x:address
	wire         mm_interconnect_0_floor2_x_s1_write;                          // mm_interconnect_0:floor2_x_s1_write -> floor2_x:write_n
	wire  [31:0] mm_interconnect_0_floor2_x_s1_writedata;                      // mm_interconnect_0:floor2_x_s1_writedata -> floor2_x:writedata
	wire         mm_interconnect_0_floor3_x_s1_chipselect;                     // mm_interconnect_0:floor3_x_s1_chipselect -> floor3_x:chipselect
	wire  [31:0] mm_interconnect_0_floor3_x_s1_readdata;                       // floor3_x:readdata -> mm_interconnect_0:floor3_x_s1_readdata
	wire   [1:0] mm_interconnect_0_floor3_x_s1_address;                        // mm_interconnect_0:floor3_x_s1_address -> floor3_x:address
	wire         mm_interconnect_0_floor3_x_s1_write;                          // mm_interconnect_0:floor3_x_s1_write -> floor3_x:write_n
	wire  [31:0] mm_interconnect_0_floor3_x_s1_writedata;                      // mm_interconnect_0:floor3_x_s1_writedata -> floor3_x:writedata
	wire         mm_interconnect_0_floor4_x_s1_chipselect;                     // mm_interconnect_0:floor4_x_s1_chipselect -> floor4_x:chipselect
	wire  [31:0] mm_interconnect_0_floor4_x_s1_readdata;                       // floor4_x:readdata -> mm_interconnect_0:floor4_x_s1_readdata
	wire   [1:0] mm_interconnect_0_floor4_x_s1_address;                        // mm_interconnect_0:floor4_x_s1_address -> floor4_x:address
	wire         mm_interconnect_0_floor4_x_s1_write;                          // mm_interconnect_0:floor4_x_s1_write -> floor4_x:write_n
	wire  [31:0] mm_interconnect_0_floor4_x_s1_writedata;                      // mm_interconnect_0:floor4_x_s1_writedata -> floor4_x:writedata
	wire         mm_interconnect_0_floor5_x_s1_chipselect;                     // mm_interconnect_0:floor5_x_s1_chipselect -> floor5_x:chipselect
	wire  [31:0] mm_interconnect_0_floor5_x_s1_readdata;                       // floor5_x:readdata -> mm_interconnect_0:floor5_x_s1_readdata
	wire   [1:0] mm_interconnect_0_floor5_x_s1_address;                        // mm_interconnect_0:floor5_x_s1_address -> floor5_x:address
	wire         mm_interconnect_0_floor5_x_s1_write;                          // mm_interconnect_0:floor5_x_s1_write -> floor5_x:write_n
	wire  [31:0] mm_interconnect_0_floor5_x_s1_writedata;                      // mm_interconnect_0:floor5_x_s1_writedata -> floor5_x:writedata
	wire         mm_interconnect_0_floor6_x_s1_chipselect;                     // mm_interconnect_0:floor6_x_s1_chipselect -> floor6_x:chipselect
	wire  [31:0] mm_interconnect_0_floor6_x_s1_readdata;                       // floor6_x:readdata -> mm_interconnect_0:floor6_x_s1_readdata
	wire   [1:0] mm_interconnect_0_floor6_x_s1_address;                        // mm_interconnect_0:floor6_x_s1_address -> floor6_x:address
	wire         mm_interconnect_0_floor6_x_s1_write;                          // mm_interconnect_0:floor6_x_s1_write -> floor6_x:write_n
	wire  [31:0] mm_interconnect_0_floor6_x_s1_writedata;                      // mm_interconnect_0:floor6_x_s1_writedata -> floor6_x:writedata
	wire         mm_interconnect_0_floor7_x_s1_chipselect;                     // mm_interconnect_0:floor7_x_s1_chipselect -> floor7_x:chipselect
	wire  [31:0] mm_interconnect_0_floor7_x_s1_readdata;                       // floor7_x:readdata -> mm_interconnect_0:floor7_x_s1_readdata
	wire   [1:0] mm_interconnect_0_floor7_x_s1_address;                        // mm_interconnect_0:floor7_x_s1_address -> floor7_x:address
	wire         mm_interconnect_0_floor7_x_s1_write;                          // mm_interconnect_0:floor7_x_s1_write -> floor7_x:write_n
	wire  [31:0] mm_interconnect_0_floor7_x_s1_writedata;                      // mm_interconnect_0:floor7_x_s1_writedata -> floor7_x:writedata
	wire         mm_interconnect_0_floor8_x_s1_chipselect;                     // mm_interconnect_0:floor8_x_s1_chipselect -> floor8_x:chipselect
	wire  [31:0] mm_interconnect_0_floor8_x_s1_readdata;                       // floor8_x:readdata -> mm_interconnect_0:floor8_x_s1_readdata
	wire   [1:0] mm_interconnect_0_floor8_x_s1_address;                        // mm_interconnect_0:floor8_x_s1_address -> floor8_x:address
	wire         mm_interconnect_0_floor8_x_s1_write;                          // mm_interconnect_0:floor8_x_s1_write -> floor8_x:write_n
	wire  [31:0] mm_interconnect_0_floor8_x_s1_writedata;                      // mm_interconnect_0:floor8_x_s1_writedata -> floor8_x:writedata
	wire         mm_interconnect_0_floor2_y_s1_chipselect;                     // mm_interconnect_0:floor2_y_s1_chipselect -> floor2_y:chipselect
	wire  [31:0] mm_interconnect_0_floor2_y_s1_readdata;                       // floor2_y:readdata -> mm_interconnect_0:floor2_y_s1_readdata
	wire   [1:0] mm_interconnect_0_floor2_y_s1_address;                        // mm_interconnect_0:floor2_y_s1_address -> floor2_y:address
	wire         mm_interconnect_0_floor2_y_s1_write;                          // mm_interconnect_0:floor2_y_s1_write -> floor2_y:write_n
	wire  [31:0] mm_interconnect_0_floor2_y_s1_writedata;                      // mm_interconnect_0:floor2_y_s1_writedata -> floor2_y:writedata
	wire         mm_interconnect_0_floor3_y_s1_chipselect;                     // mm_interconnect_0:floor3_y_s1_chipselect -> floor3_y:chipselect
	wire  [31:0] mm_interconnect_0_floor3_y_s1_readdata;                       // floor3_y:readdata -> mm_interconnect_0:floor3_y_s1_readdata
	wire   [1:0] mm_interconnect_0_floor3_y_s1_address;                        // mm_interconnect_0:floor3_y_s1_address -> floor3_y:address
	wire         mm_interconnect_0_floor3_y_s1_write;                          // mm_interconnect_0:floor3_y_s1_write -> floor3_y:write_n
	wire  [31:0] mm_interconnect_0_floor3_y_s1_writedata;                      // mm_interconnect_0:floor3_y_s1_writedata -> floor3_y:writedata
	wire         mm_interconnect_0_floor4_y_s1_chipselect;                     // mm_interconnect_0:floor4_y_s1_chipselect -> floor4_y:chipselect
	wire  [31:0] mm_interconnect_0_floor4_y_s1_readdata;                       // floor4_y:readdata -> mm_interconnect_0:floor4_y_s1_readdata
	wire   [1:0] mm_interconnect_0_floor4_y_s1_address;                        // mm_interconnect_0:floor4_y_s1_address -> floor4_y:address
	wire         mm_interconnect_0_floor4_y_s1_write;                          // mm_interconnect_0:floor4_y_s1_write -> floor4_y:write_n
	wire  [31:0] mm_interconnect_0_floor4_y_s1_writedata;                      // mm_interconnect_0:floor4_y_s1_writedata -> floor4_y:writedata
	wire         mm_interconnect_0_floor5_y_s1_chipselect;                     // mm_interconnect_0:floor5_y_s1_chipselect -> floor5_y:chipselect
	wire  [31:0] mm_interconnect_0_floor5_y_s1_readdata;                       // floor5_y:readdata -> mm_interconnect_0:floor5_y_s1_readdata
	wire   [1:0] mm_interconnect_0_floor5_y_s1_address;                        // mm_interconnect_0:floor5_y_s1_address -> floor5_y:address
	wire         mm_interconnect_0_floor5_y_s1_write;                          // mm_interconnect_0:floor5_y_s1_write -> floor5_y:write_n
	wire  [31:0] mm_interconnect_0_floor5_y_s1_writedata;                      // mm_interconnect_0:floor5_y_s1_writedata -> floor5_y:writedata
	wire         mm_interconnect_0_floor6_y_s1_chipselect;                     // mm_interconnect_0:floor6_y_s1_chipselect -> floor6_y:chipselect
	wire  [31:0] mm_interconnect_0_floor6_y_s1_readdata;                       // floor6_y:readdata -> mm_interconnect_0:floor6_y_s1_readdata
	wire   [1:0] mm_interconnect_0_floor6_y_s1_address;                        // mm_interconnect_0:floor6_y_s1_address -> floor6_y:address
	wire         mm_interconnect_0_floor6_y_s1_write;                          // mm_interconnect_0:floor6_y_s1_write -> floor6_y:write_n
	wire  [31:0] mm_interconnect_0_floor6_y_s1_writedata;                      // mm_interconnect_0:floor6_y_s1_writedata -> floor6_y:writedata
	wire         mm_interconnect_0_floor7_y_s1_chipselect;                     // mm_interconnect_0:floor7_y_s1_chipselect -> floor7_y:chipselect
	wire  [31:0] mm_interconnect_0_floor7_y_s1_readdata;                       // floor7_y:readdata -> mm_interconnect_0:floor7_y_s1_readdata
	wire   [1:0] mm_interconnect_0_floor7_y_s1_address;                        // mm_interconnect_0:floor7_y_s1_address -> floor7_y:address
	wire         mm_interconnect_0_floor7_y_s1_write;                          // mm_interconnect_0:floor7_y_s1_write -> floor7_y:write_n
	wire  [31:0] mm_interconnect_0_floor7_y_s1_writedata;                      // mm_interconnect_0:floor7_y_s1_writedata -> floor7_y:writedata
	wire         mm_interconnect_0_floor8_y_s1_chipselect;                     // mm_interconnect_0:floor8_y_s1_chipselect -> floor8_y:chipselect
	wire  [31:0] mm_interconnect_0_floor8_y_s1_readdata;                       // floor8_y:readdata -> mm_interconnect_0:floor8_y_s1_readdata
	wire   [1:0] mm_interconnect_0_floor8_y_s1_address;                        // mm_interconnect_0:floor8_y_s1_address -> floor8_y:address
	wire         mm_interconnect_0_floor8_y_s1_write;                          // mm_interconnect_0:floor8_y_s1_write -> floor8_y:write_n
	wire  [31:0] mm_interconnect_0_floor8_y_s1_writedata;                      // mm_interconnect_0:floor8_y_s1_writedata -> floor8_y:writedata
	wire         mm_interconnect_0_score_s1_chipselect;                        // mm_interconnect_0:score_s1_chipselect -> score:chipselect
	wire  [31:0] mm_interconnect_0_score_s1_readdata;                          // score:readdata -> mm_interconnect_0:score_s1_readdata
	wire   [1:0] mm_interconnect_0_score_s1_address;                           // mm_interconnect_0:score_s1_address -> score:address
	wire         mm_interconnect_0_score_s1_write;                             // mm_interconnect_0:score_s1_write -> score:write_n
	wire  [31:0] mm_interconnect_0_score_s1_writedata;                         // mm_interconnect_0:score_s1_writedata -> score:writedata
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [doodle_x:reset_n, doodle_y:reset_n, floor1_x:reset_n, floor1_y:reset_n, floor2_x:reset_n, floor2_y:reset_n, floor3_x:reset_n, floor3_y:reset_n, floor4_x:reset_n, floor4_y:reset_n, floor5_x:reset_n, floor5_y:reset_n, floor6_x:reset_n, floor6_y:reset_n, floor7_x:reset_n, floor7_y:reset_n, floor8_x:reset_n, floor8_y:reset_n, jtag_uart_0:rst_n, keycode:reset_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, otg_hpi_address:reset_n, otg_hpi_cs:reset_n, otg_hpi_data:reset_n, otg_hpi_r:reset_n, otg_hpi_reset:reset_n, otg_hpi_w:reset_n, score:reset_n]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram_pll:reset, sysid_qsys_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                       // rst_controller_001:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                           // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	nios_system_doodle_x doodle_x (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_doodle_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_doodle_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_doodle_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_doodle_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_doodle_x_s1_readdata),   //                    .readdata
		.out_port   (doodle_x_export)                           // external_connection.export
	);

	nios_system_doodle_x doodle_y (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_doodle_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_doodle_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_doodle_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_doodle_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_doodle_y_s1_readdata),   //                    .readdata
		.out_port   (doodle_y_export)                           // external_connection.export
	);

	nios_system_doodle_x floor1_x (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor1_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor1_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor1_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor1_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor1_x_s1_readdata),   //                    .readdata
		.out_port   (floor1_x_export)                           // external_connection.export
	);

	nios_system_doodle_x floor1_y (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor1_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor1_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor1_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor1_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor1_y_s1_readdata),   //                    .readdata
		.out_port   (floor1_y_export)                           // external_connection.export
	);

	nios_system_doodle_x floor2_x (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor2_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor2_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor2_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor2_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor2_x_s1_readdata),   //                    .readdata
		.out_port   (floor2_x_export)                           // external_connection.export
	);

	nios_system_doodle_x floor2_y (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor2_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor2_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor2_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor2_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor2_y_s1_readdata),   //                    .readdata
		.out_port   (floor2_y_export)                           // external_connection.export
	);

	nios_system_doodle_x floor3_x (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor3_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor3_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor3_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor3_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor3_x_s1_readdata),   //                    .readdata
		.out_port   (floor3_x_export)                           // external_connection.export
	);

	nios_system_doodle_x floor3_y (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor3_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor3_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor3_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor3_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor3_y_s1_readdata),   //                    .readdata
		.out_port   (floor3_y_export)                           // external_connection.export
	);

	nios_system_doodle_x floor4_x (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor4_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor4_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor4_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor4_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor4_x_s1_readdata),   //                    .readdata
		.out_port   (floor4_x_export)                           // external_connection.export
	);

	nios_system_doodle_x floor4_y (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor4_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor4_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor4_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor4_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor4_y_s1_readdata),   //                    .readdata
		.out_port   (floor4_y_export)                           // external_connection.export
	);

	nios_system_doodle_x floor5_x (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor5_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor5_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor5_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor5_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor5_x_s1_readdata),   //                    .readdata
		.out_port   (floor5_x_export)                           // external_connection.export
	);

	nios_system_doodle_x floor5_y (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor5_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor5_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor5_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor5_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor5_y_s1_readdata),   //                    .readdata
		.out_port   (floor5_y_export)                           // external_connection.export
	);

	nios_system_doodle_x floor6_x (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor6_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor6_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor6_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor6_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor6_x_s1_readdata),   //                    .readdata
		.out_port   (floor6_x_export)                           // external_connection.export
	);

	nios_system_doodle_x floor6_y (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor6_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor6_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor6_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor6_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor6_y_s1_readdata),   //                    .readdata
		.out_port   (floor6_y_export)                           // external_connection.export
	);

	nios_system_doodle_x floor7_x (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor7_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor7_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor7_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor7_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor7_x_s1_readdata),   //                    .readdata
		.out_port   (floor7_x_export)                           // external_connection.export
	);

	nios_system_doodle_x floor7_y (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor7_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor7_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor7_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor7_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor7_y_s1_readdata),   //                    .readdata
		.out_port   (floor7_y_export)                           // external_connection.export
	);

	nios_system_doodle_x floor8_x (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor8_x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor8_x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor8_x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor8_x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor8_x_s1_readdata),   //                    .readdata
		.out_port   (floor8_x_export)                           // external_connection.export
	);

	nios_system_doodle_x floor8_y (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_floor8_y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_floor8_y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_floor8_y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_floor8_y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_floor8_y_s1_readdata),   //                    .readdata
		.out_port   (floor8_y_export)                           // external_connection.export
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_keycode keycode (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_keycode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_s1_readdata),   //                    .readdata
		.out_port   (keycode_export)                           // external_connection.export
	);

	nios_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                          //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),                       //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios_system_otg_hpi_address otg_hpi_address (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	nios_system_otg_hpi_cs otg_hpi_cs (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	nios_system_otg_hpi_data otg_hpi_data (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	nios_system_otg_hpi_cs otg_hpi_r (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	nios_system_otg_hpi_cs otg_hpi_reset (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_reset_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_reset_export)                           // external_connection.export
	);

	nios_system_otg_hpi_cs otg_hpi_w (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	nios_system_score score (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_score_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_score_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_score_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_score_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_score_s1_readdata),   //                    .readdata
		.out_port   (score_export)                           // external_connection.export
	);

	nios_system_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	nios_system_sdram_pll sdram_pll (
		.clk                (clk_clk),                                         //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),              // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                                   //                    c1.clk
		.scandone           (),                                                //           (terminated)
		.scandataout        (),                                                //           (terminated)
		.areset             (1'b0),                                            //           (terminated)
		.locked             (),                                                //           (terminated)
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (4'b0000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0),                                            //           (terminated)
		.scanclkena         (1'b0),                                            //           (terminated)
		.scandata           (1'b0),                                            //           (terminated)
		.configupdate       (1'b0)                                             //           (terminated)
	);

	nios_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.sdram_pll_c0_clk                                 (sdram_pll_c0_clk),                                             //                               sdram_pll_c0.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                               //    jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                           // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset          (rst_controller_002_reset_out_reset),                           //          sdram_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.doodle_x_s1_address                              (mm_interconnect_0_doodle_x_s1_address),                        //                                doodle_x_s1.address
		.doodle_x_s1_write                                (mm_interconnect_0_doodle_x_s1_write),                          //                                           .write
		.doodle_x_s1_readdata                             (mm_interconnect_0_doodle_x_s1_readdata),                       //                                           .readdata
		.doodle_x_s1_writedata                            (mm_interconnect_0_doodle_x_s1_writedata),                      //                                           .writedata
		.doodle_x_s1_chipselect                           (mm_interconnect_0_doodle_x_s1_chipselect),                     //                                           .chipselect
		.doodle_y_s1_address                              (mm_interconnect_0_doodle_y_s1_address),                        //                                doodle_y_s1.address
		.doodle_y_s1_write                                (mm_interconnect_0_doodle_y_s1_write),                          //                                           .write
		.doodle_y_s1_readdata                             (mm_interconnect_0_doodle_y_s1_readdata),                       //                                           .readdata
		.doodle_y_s1_writedata                            (mm_interconnect_0_doodle_y_s1_writedata),                      //                                           .writedata
		.doodle_y_s1_chipselect                           (mm_interconnect_0_doodle_y_s1_chipselect),                     //                                           .chipselect
		.floor1_x_s1_address                              (mm_interconnect_0_floor1_x_s1_address),                        //                                floor1_x_s1.address
		.floor1_x_s1_write                                (mm_interconnect_0_floor1_x_s1_write),                          //                                           .write
		.floor1_x_s1_readdata                             (mm_interconnect_0_floor1_x_s1_readdata),                       //                                           .readdata
		.floor1_x_s1_writedata                            (mm_interconnect_0_floor1_x_s1_writedata),                      //                                           .writedata
		.floor1_x_s1_chipselect                           (mm_interconnect_0_floor1_x_s1_chipselect),                     //                                           .chipselect
		.floor1_y_s1_address                              (mm_interconnect_0_floor1_y_s1_address),                        //                                floor1_y_s1.address
		.floor1_y_s1_write                                (mm_interconnect_0_floor1_y_s1_write),                          //                                           .write
		.floor1_y_s1_readdata                             (mm_interconnect_0_floor1_y_s1_readdata),                       //                                           .readdata
		.floor1_y_s1_writedata                            (mm_interconnect_0_floor1_y_s1_writedata),                      //                                           .writedata
		.floor1_y_s1_chipselect                           (mm_interconnect_0_floor1_y_s1_chipselect),                     //                                           .chipselect
		.floor2_x_s1_address                              (mm_interconnect_0_floor2_x_s1_address),                        //                                floor2_x_s1.address
		.floor2_x_s1_write                                (mm_interconnect_0_floor2_x_s1_write),                          //                                           .write
		.floor2_x_s1_readdata                             (mm_interconnect_0_floor2_x_s1_readdata),                       //                                           .readdata
		.floor2_x_s1_writedata                            (mm_interconnect_0_floor2_x_s1_writedata),                      //                                           .writedata
		.floor2_x_s1_chipselect                           (mm_interconnect_0_floor2_x_s1_chipselect),                     //                                           .chipselect
		.floor2_y_s1_address                              (mm_interconnect_0_floor2_y_s1_address),                        //                                floor2_y_s1.address
		.floor2_y_s1_write                                (mm_interconnect_0_floor2_y_s1_write),                          //                                           .write
		.floor2_y_s1_readdata                             (mm_interconnect_0_floor2_y_s1_readdata),                       //                                           .readdata
		.floor2_y_s1_writedata                            (mm_interconnect_0_floor2_y_s1_writedata),                      //                                           .writedata
		.floor2_y_s1_chipselect                           (mm_interconnect_0_floor2_y_s1_chipselect),                     //                                           .chipselect
		.floor3_x_s1_address                              (mm_interconnect_0_floor3_x_s1_address),                        //                                floor3_x_s1.address
		.floor3_x_s1_write                                (mm_interconnect_0_floor3_x_s1_write),                          //                                           .write
		.floor3_x_s1_readdata                             (mm_interconnect_0_floor3_x_s1_readdata),                       //                                           .readdata
		.floor3_x_s1_writedata                            (mm_interconnect_0_floor3_x_s1_writedata),                      //                                           .writedata
		.floor3_x_s1_chipselect                           (mm_interconnect_0_floor3_x_s1_chipselect),                     //                                           .chipselect
		.floor3_y_s1_address                              (mm_interconnect_0_floor3_y_s1_address),                        //                                floor3_y_s1.address
		.floor3_y_s1_write                                (mm_interconnect_0_floor3_y_s1_write),                          //                                           .write
		.floor3_y_s1_readdata                             (mm_interconnect_0_floor3_y_s1_readdata),                       //                                           .readdata
		.floor3_y_s1_writedata                            (mm_interconnect_0_floor3_y_s1_writedata),                      //                                           .writedata
		.floor3_y_s1_chipselect                           (mm_interconnect_0_floor3_y_s1_chipselect),                     //                                           .chipselect
		.floor4_x_s1_address                              (mm_interconnect_0_floor4_x_s1_address),                        //                                floor4_x_s1.address
		.floor4_x_s1_write                                (mm_interconnect_0_floor4_x_s1_write),                          //                                           .write
		.floor4_x_s1_readdata                             (mm_interconnect_0_floor4_x_s1_readdata),                       //                                           .readdata
		.floor4_x_s1_writedata                            (mm_interconnect_0_floor4_x_s1_writedata),                      //                                           .writedata
		.floor4_x_s1_chipselect                           (mm_interconnect_0_floor4_x_s1_chipselect),                     //                                           .chipselect
		.floor4_y_s1_address                              (mm_interconnect_0_floor4_y_s1_address),                        //                                floor4_y_s1.address
		.floor4_y_s1_write                                (mm_interconnect_0_floor4_y_s1_write),                          //                                           .write
		.floor4_y_s1_readdata                             (mm_interconnect_0_floor4_y_s1_readdata),                       //                                           .readdata
		.floor4_y_s1_writedata                            (mm_interconnect_0_floor4_y_s1_writedata),                      //                                           .writedata
		.floor4_y_s1_chipselect                           (mm_interconnect_0_floor4_y_s1_chipselect),                     //                                           .chipselect
		.floor5_x_s1_address                              (mm_interconnect_0_floor5_x_s1_address),                        //                                floor5_x_s1.address
		.floor5_x_s1_write                                (mm_interconnect_0_floor5_x_s1_write),                          //                                           .write
		.floor5_x_s1_readdata                             (mm_interconnect_0_floor5_x_s1_readdata),                       //                                           .readdata
		.floor5_x_s1_writedata                            (mm_interconnect_0_floor5_x_s1_writedata),                      //                                           .writedata
		.floor5_x_s1_chipselect                           (mm_interconnect_0_floor5_x_s1_chipselect),                     //                                           .chipselect
		.floor5_y_s1_address                              (mm_interconnect_0_floor5_y_s1_address),                        //                                floor5_y_s1.address
		.floor5_y_s1_write                                (mm_interconnect_0_floor5_y_s1_write),                          //                                           .write
		.floor5_y_s1_readdata                             (mm_interconnect_0_floor5_y_s1_readdata),                       //                                           .readdata
		.floor5_y_s1_writedata                            (mm_interconnect_0_floor5_y_s1_writedata),                      //                                           .writedata
		.floor5_y_s1_chipselect                           (mm_interconnect_0_floor5_y_s1_chipselect),                     //                                           .chipselect
		.floor6_x_s1_address                              (mm_interconnect_0_floor6_x_s1_address),                        //                                floor6_x_s1.address
		.floor6_x_s1_write                                (mm_interconnect_0_floor6_x_s1_write),                          //                                           .write
		.floor6_x_s1_readdata                             (mm_interconnect_0_floor6_x_s1_readdata),                       //                                           .readdata
		.floor6_x_s1_writedata                            (mm_interconnect_0_floor6_x_s1_writedata),                      //                                           .writedata
		.floor6_x_s1_chipselect                           (mm_interconnect_0_floor6_x_s1_chipselect),                     //                                           .chipselect
		.floor6_y_s1_address                              (mm_interconnect_0_floor6_y_s1_address),                        //                                floor6_y_s1.address
		.floor6_y_s1_write                                (mm_interconnect_0_floor6_y_s1_write),                          //                                           .write
		.floor6_y_s1_readdata                             (mm_interconnect_0_floor6_y_s1_readdata),                       //                                           .readdata
		.floor6_y_s1_writedata                            (mm_interconnect_0_floor6_y_s1_writedata),                      //                                           .writedata
		.floor6_y_s1_chipselect                           (mm_interconnect_0_floor6_y_s1_chipselect),                     //                                           .chipselect
		.floor7_x_s1_address                              (mm_interconnect_0_floor7_x_s1_address),                        //                                floor7_x_s1.address
		.floor7_x_s1_write                                (mm_interconnect_0_floor7_x_s1_write),                          //                                           .write
		.floor7_x_s1_readdata                             (mm_interconnect_0_floor7_x_s1_readdata),                       //                                           .readdata
		.floor7_x_s1_writedata                            (mm_interconnect_0_floor7_x_s1_writedata),                      //                                           .writedata
		.floor7_x_s1_chipselect                           (mm_interconnect_0_floor7_x_s1_chipselect),                     //                                           .chipselect
		.floor7_y_s1_address                              (mm_interconnect_0_floor7_y_s1_address),                        //                                floor7_y_s1.address
		.floor7_y_s1_write                                (mm_interconnect_0_floor7_y_s1_write),                          //                                           .write
		.floor7_y_s1_readdata                             (mm_interconnect_0_floor7_y_s1_readdata),                       //                                           .readdata
		.floor7_y_s1_writedata                            (mm_interconnect_0_floor7_y_s1_writedata),                      //                                           .writedata
		.floor7_y_s1_chipselect                           (mm_interconnect_0_floor7_y_s1_chipselect),                     //                                           .chipselect
		.floor8_x_s1_address                              (mm_interconnect_0_floor8_x_s1_address),                        //                                floor8_x_s1.address
		.floor8_x_s1_write                                (mm_interconnect_0_floor8_x_s1_write),                          //                                           .write
		.floor8_x_s1_readdata                             (mm_interconnect_0_floor8_x_s1_readdata),                       //                                           .readdata
		.floor8_x_s1_writedata                            (mm_interconnect_0_floor8_x_s1_writedata),                      //                                           .writedata
		.floor8_x_s1_chipselect                           (mm_interconnect_0_floor8_x_s1_chipselect),                     //                                           .chipselect
		.floor8_y_s1_address                              (mm_interconnect_0_floor8_y_s1_address),                        //                                floor8_y_s1.address
		.floor8_y_s1_write                                (mm_interconnect_0_floor8_y_s1_write),                          //                                           .write
		.floor8_y_s1_readdata                             (mm_interconnect_0_floor8_y_s1_readdata),                       //                                           .readdata
		.floor8_y_s1_writedata                            (mm_interconnect_0_floor8_y_s1_writedata),                      //                                           .writedata
		.floor8_y_s1_chipselect                           (mm_interconnect_0_floor8_y_s1_chipselect),                     //                                           .chipselect
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.keycode_s1_address                               (mm_interconnect_0_keycode_s1_address),                         //                                 keycode_s1.address
		.keycode_s1_write                                 (mm_interconnect_0_keycode_s1_write),                           //                                           .write
		.keycode_s1_readdata                              (mm_interconnect_0_keycode_s1_readdata),                        //                                           .readdata
		.keycode_s1_writedata                             (mm_interconnect_0_keycode_s1_writedata),                       //                                           .writedata
		.keycode_s1_chipselect                            (mm_interconnect_0_keycode_s1_chipselect),                      //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                  //                                           .clken
		.otg_hpi_address_s1_address                       (mm_interconnect_0_otg_hpi_address_s1_address),                 //                         otg_hpi_address_s1.address
		.otg_hpi_address_s1_write                         (mm_interconnect_0_otg_hpi_address_s1_write),                   //                                           .write
		.otg_hpi_address_s1_readdata                      (mm_interconnect_0_otg_hpi_address_s1_readdata),                //                                           .readdata
		.otg_hpi_address_s1_writedata                     (mm_interconnect_0_otg_hpi_address_s1_writedata),               //                                           .writedata
		.otg_hpi_address_s1_chipselect                    (mm_interconnect_0_otg_hpi_address_s1_chipselect),              //                                           .chipselect
		.otg_hpi_cs_s1_address                            (mm_interconnect_0_otg_hpi_cs_s1_address),                      //                              otg_hpi_cs_s1.address
		.otg_hpi_cs_s1_write                              (mm_interconnect_0_otg_hpi_cs_s1_write),                        //                                           .write
		.otg_hpi_cs_s1_readdata                           (mm_interconnect_0_otg_hpi_cs_s1_readdata),                     //                                           .readdata
		.otg_hpi_cs_s1_writedata                          (mm_interconnect_0_otg_hpi_cs_s1_writedata),                    //                                           .writedata
		.otg_hpi_cs_s1_chipselect                         (mm_interconnect_0_otg_hpi_cs_s1_chipselect),                   //                                           .chipselect
		.otg_hpi_data_s1_address                          (mm_interconnect_0_otg_hpi_data_s1_address),                    //                            otg_hpi_data_s1.address
		.otg_hpi_data_s1_write                            (mm_interconnect_0_otg_hpi_data_s1_write),                      //                                           .write
		.otg_hpi_data_s1_readdata                         (mm_interconnect_0_otg_hpi_data_s1_readdata),                   //                                           .readdata
		.otg_hpi_data_s1_writedata                        (mm_interconnect_0_otg_hpi_data_s1_writedata),                  //                                           .writedata
		.otg_hpi_data_s1_chipselect                       (mm_interconnect_0_otg_hpi_data_s1_chipselect),                 //                                           .chipselect
		.otg_hpi_r_s1_address                             (mm_interconnect_0_otg_hpi_r_s1_address),                       //                               otg_hpi_r_s1.address
		.otg_hpi_r_s1_write                               (mm_interconnect_0_otg_hpi_r_s1_write),                         //                                           .write
		.otg_hpi_r_s1_readdata                            (mm_interconnect_0_otg_hpi_r_s1_readdata),                      //                                           .readdata
		.otg_hpi_r_s1_writedata                           (mm_interconnect_0_otg_hpi_r_s1_writedata),                     //                                           .writedata
		.otg_hpi_r_s1_chipselect                          (mm_interconnect_0_otg_hpi_r_s1_chipselect),                    //                                           .chipselect
		.otg_hpi_reset_s1_address                         (mm_interconnect_0_otg_hpi_reset_s1_address),                   //                           otg_hpi_reset_s1.address
		.otg_hpi_reset_s1_write                           (mm_interconnect_0_otg_hpi_reset_s1_write),                     //                                           .write
		.otg_hpi_reset_s1_readdata                        (mm_interconnect_0_otg_hpi_reset_s1_readdata),                  //                                           .readdata
		.otg_hpi_reset_s1_writedata                       (mm_interconnect_0_otg_hpi_reset_s1_writedata),                 //                                           .writedata
		.otg_hpi_reset_s1_chipselect                      (mm_interconnect_0_otg_hpi_reset_s1_chipselect),                //                                           .chipselect
		.otg_hpi_w_s1_address                             (mm_interconnect_0_otg_hpi_w_s1_address),                       //                               otg_hpi_w_s1.address
		.otg_hpi_w_s1_write                               (mm_interconnect_0_otg_hpi_w_s1_write),                         //                                           .write
		.otg_hpi_w_s1_readdata                            (mm_interconnect_0_otg_hpi_w_s1_readdata),                      //                                           .readdata
		.otg_hpi_w_s1_writedata                           (mm_interconnect_0_otg_hpi_w_s1_writedata),                     //                                           .writedata
		.otg_hpi_w_s1_chipselect                          (mm_interconnect_0_otg_hpi_w_s1_chipselect),                    //                                           .chipselect
		.score_s1_address                                 (mm_interconnect_0_score_s1_address),                           //                                   score_s1.address
		.score_s1_write                                   (mm_interconnect_0_score_s1_write),                             //                                           .write
		.score_s1_readdata                                (mm_interconnect_0_score_s1_readdata),                          //                                           .readdata
		.score_s1_writedata                               (mm_interconnect_0_score_s1_writedata),                         //                                           .writedata
		.score_s1_chipselect                              (mm_interconnect_0_score_s1_chipselect),                        //                                           .chipselect
		.sdram_s1_address                                 (mm_interconnect_0_sdram_s1_address),                           //                                   sdram_s1.address
		.sdram_s1_write                                   (mm_interconnect_0_sdram_s1_write),                             //                                           .write
		.sdram_s1_read                                    (mm_interconnect_0_sdram_s1_read),                              //                                           .read
		.sdram_s1_readdata                                (mm_interconnect_0_sdram_s1_readdata),                          //                                           .readdata
		.sdram_s1_writedata                               (mm_interconnect_0_sdram_s1_writedata),                         //                                           .writedata
		.sdram_s1_byteenable                              (mm_interconnect_0_sdram_s1_byteenable),                        //                                           .byteenable
		.sdram_s1_readdatavalid                           (mm_interconnect_0_sdram_s1_readdatavalid),                     //                                           .readdatavalid
		.sdram_s1_waitrequest                             (mm_interconnect_0_sdram_s1_waitrequest),                       //                                           .waitrequest
		.sdram_s1_chipselect                              (mm_interconnect_0_sdram_s1_chipselect),                        //                                           .chipselect
		.sdram_pll_pll_slave_address                      (mm_interconnect_0_sdram_pll_pll_slave_address),                //                        sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                        (mm_interconnect_0_sdram_pll_pll_slave_write),                  //                                           .write
		.sdram_pll_pll_slave_read                         (mm_interconnect_0_sdram_pll_pll_slave_read),                   //                                           .read
		.sdram_pll_pll_slave_readdata                     (mm_interconnect_0_sdram_pll_pll_slave_readdata),               //                                           .readdata
		.sdram_pll_pll_slave_writedata                    (mm_interconnect_0_sdram_pll_pll_slave_writedata),              //                                           .writedata
		.sysid_qsys_0_control_slave_address               (mm_interconnect_0_sysid_qsys_0_control_slave_address),         //                 sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata              (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)         //                                           .readdata
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (sdram_pll_c0_clk),                           //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
